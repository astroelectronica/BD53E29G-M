.title KiCad schematic
.include "C:/AE/BD53E29G/models/BD53E29G.lib"
.include "C:/AE/BD53E29G/models/C2012C0G2W101J060AA_p.mod"
.include "C:/AE/BD53E29G/models/C2012JB2E102M085AA_p.mod"
.include "C:/AE/BD53E29G/models/C2012X7R2A104M125AA_p.mod"
XU4 /OUT 0 C2012JB2E102M085AA_p
XU1 /OUT VDD 0 unconnected-_U1-PadNC_ /CT BD53E29G
V1 VDD 0 {VSUPPLY}
XU3 /CT 0 C2012C0G2W101J060AA_p
XU2 VDD 0 C2012X7R2A104M125AA_p
.end
